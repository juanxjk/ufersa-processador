LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY processador IS
	PORT(
		clk, rst			: IN STD_LOGIC;
	);
END ENTITY;

ARCHITECTURE comportamento OF processador IS
COMPONENT -- !!!!!!!!!!!!!!!!!!!!!!!!!

END COMPONENT;

COMPONENT -- !!!!!!!!!!!!!!!!!!!!!!!!!

END COMPONENT;

COMPONENT -- !!!!!!!!!!!!!!!!!!!!!!!!!

END COMPONENT;

SIGNAL -- !!!!!!!!!!!!!!!!!!!!!!!!!

BEGIN 
	
	port map() -- !!!!!!!!!!!!!!!!!!!!!!!!!
END comportamento;